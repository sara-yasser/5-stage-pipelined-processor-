LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE ieee.numeric_std.all; 

entity compare_logic is
port
(
    

    );
end entity;

architecture compare_logic_arc of compare_logic is

    begin
        
end architecture;

